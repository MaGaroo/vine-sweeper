module Receiver #(parameter clockperbit) (rxdata, rxfinish, rx, clock, reset);
	input clock, reset, rx;
	output reg rxfinish;
	output reg [7:0] rxdata;
	
	

endmodule
