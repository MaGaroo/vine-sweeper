module minesweeper(out, in);
	output out;
	input in;

	
	
endmodule
