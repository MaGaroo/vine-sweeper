module Receiver #(parameter clockperbit) (rxdata, rxfinish, rx, clock, reset);
	

endmodule
